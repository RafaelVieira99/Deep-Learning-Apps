-- DE2_115_SD_CARD_NIOS.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE2_115_SD_CARD_NIOS is
	port (
		activations_index_external_connection_export                    : out   std_logic_vector(3 downto 0);                     --     activations_index_external_connection.export
		altpll_areset_conduit_export                                    : in    std_logic                     := '0';             --                     altpll_areset_conduit.export
		altpll_c1_clk                                                   : out   std_logic;                                        --                                 altpll_c1.clk
		altpll_c3_clk                                                   : out   std_logic;                                        --                                 altpll_c3.clk
		altpll_locked_conduit_export                                    : out   std_logic;                                        --                     altpll_locked_conduit.export
		c0_out_clk_clk                                                  : out   std_logic;                                        --                                c0_out_clk.clk
		c2_out_clk_clk                                                  : out   std_logic;                                        --                                c2_out_clk.clk
		clk_50_clk_in_clk                                               : in    std_logic                     := '0';             --                             clk_50_clk_in.clk
		floatdata_output_external_connection_export                     : out   std_logic_vector(31 downto 0);                    --      floatdata_output_external_connection.export
		key_external_connection_export                                  : in    std_logic_vector(3 downto 0)  := (others => '0'); --                   key_external_connection.export
		ledg_external_connection_export                                 : out   std_logic_vector(8 downto 0);                     --                  ledg_external_connection.export
		ledr_external_connection_export                                 : out   std_logic_vector(17 downto 0);                    --                  ledr_external_connection.export
		pixel_index_external_connection_export                          : out   std_logic_vector(9 downto 0);                     --           pixel_index_external_connection.export
		reset_reset_n                                                   : in    std_logic                     := '0';             --                                     reset.reset_n
		results_input_external_connection_export                        : in    std_logic_vector(31 downto 0) := (others => '0'); --         results_input_external_connection.export
		sd_clk_external_connection_export                               : out   std_logic;                                        --                sd_clk_external_connection.export
		sd_cmd_external_connection_export                               : inout std_logic                     := '0';             --                sd_cmd_external_connection.export
		sd_dat_external_connection_export                               : inout std_logic_vector(3 downto 0)  := (others => '0'); --                sd_dat_external_connection.export
		sd_wp_n_external_connection_export                              : in    std_logic                     := '0';             --               sd_wp_n_external_connection.export
		sw_external_connection_export                                   : in    std_logic_vector(17 downto 0) := (others => '0'); --                    sw_external_connection.export
		sync_data_external_connection_export                            : out   std_logic_vector(15 downto 0);                    --             sync_data_external_connection.export
		tri_state_bridge_flash_bridge_0_out_address_to_the_cfi_flash    : out   std_logic_vector(22 downto 0);                    --       tri_state_bridge_flash_bridge_0_out.address_to_the_cfi_flash
		tri_state_bridge_flash_bridge_0_out_tri_state_bridge_flash_data : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                          .tri_state_bridge_flash_data
		tri_state_bridge_flash_bridge_0_out_write_n_to_the_cfi_flash    : out   std_logic_vector(0 downto 0);                     --                                          .write_n_to_the_cfi_flash
		tri_state_bridge_flash_bridge_0_out_select_n_to_the_cfi_flash   : out   std_logic_vector(0 downto 0);                     --                                          .select_n_to_the_cfi_flash
		tri_state_bridge_flash_bridge_0_out_read_n_to_the_cfi_flash     : out   std_logic_vector(0 downto 0);                     --                                          .read_n_to_the_cfi_flash
		video_vga_controller_0_external_interface_CLK                   : out   std_logic;                                        -- video_vga_controller_0_external_interface.CLK
		video_vga_controller_0_external_interface_HS                    : out   std_logic;                                        --                                          .HS
		video_vga_controller_0_external_interface_VS                    : out   std_logic;                                        --                                          .VS
		video_vga_controller_0_external_interface_BLANK                 : out   std_logic;                                        --                                          .BLANK
		video_vga_controller_0_external_interface_SYNC                  : out   std_logic;                                        --                                          .SYNC
		video_vga_controller_0_external_interface_R                     : out   std_logic_vector(7 downto 0);                     --                                          .R
		video_vga_controller_0_external_interface_G                     : out   std_logic_vector(7 downto 0);                     --                                          .G
		video_vga_controller_0_external_interface_B                     : out   std_logic_vector(7 downto 0);                     --                                          .B
		weight_index_external_connection_export                         : out   std_logic_vector(12 downto 0)                     --          weight_index_external_connection.export
	);
end entity DE2_115_SD_CARD_NIOS;

architecture rtl of DE2_115_SD_CARD_NIOS is
	component DE2_115_SD_CARD_NIOS_activations_index is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component DE2_115_SD_CARD_NIOS_activations_index;

	component DE2_115_SD_CARD_NIOS_altpll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X';             -- export
			phasedone          : out std_logic                                         -- export
		);
	end component DE2_115_SD_CARD_NIOS_altpll;

	component DE2_115_SD_CARD_NIOS_cfi_flash is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			uas_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_read_n_out       : out std_logic;                                        -- read_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(22 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(7 downto 0);                     -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- data_in
		);
	end component DE2_115_SD_CARD_NIOS_cfi_flash;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(8 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component DE2_115_SD_CARD_NIOS_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(25 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component DE2_115_SD_CARD_NIOS_cpu;

	component DE2_115_SD_CARD_NIOS_floatdata_output is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component DE2_115_SD_CARD_NIOS_floatdata_output;

	component DE2_115_SD_CARD_NIOS_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DE2_115_SD_CARD_NIOS_jtag_uart;

	component DE2_115_SD_CARD_NIOS_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component DE2_115_SD_CARD_NIOS_key;

	component DE2_115_SD_CARD_NIOS_ledg is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component DE2_115_SD_CARD_NIOS_ledg;

	component DE2_115_SD_CARD_NIOS_ledr is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component DE2_115_SD_CARD_NIOS_ledr;

	component DE2_115_SD_CARD_NIOS_onchip_memory2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component DE2_115_SD_CARD_NIOS_onchip_memory2;

	component DE2_115_SD_CARD_NIOS_pixel_index is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component DE2_115_SD_CARD_NIOS_pixel_index;

	component DE2_115_SD_CARD_NIOS_results_input is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component DE2_115_SD_CARD_NIOS_results_input;

	component DE2_115_SD_CARD_NIOS_sd_clk is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component DE2_115_SD_CARD_NIOS_sd_clk;

	component DE2_115_SD_CARD_NIOS_sd_cmd is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component DE2_115_SD_CARD_NIOS_sd_cmd;

	component DE2_115_SD_CARD_NIOS_sd_dat is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component DE2_115_SD_CARD_NIOS_sd_dat;

	component DE2_115_SD_CARD_NIOS_sd_wp_n is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component DE2_115_SD_CARD_NIOS_sd_wp_n;

	component DE2_115_SD_CARD_NIOS_sw is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(17 downto 0) := (others => 'X')  -- export
		);
	end component DE2_115_SD_CARD_NIOS_sw;

	component DE2_115_SD_CARD_NIOS_sync_data is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component DE2_115_SD_CARD_NIOS_sync_data;

	component DE2_115_SD_CARD_NIOS_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DE2_115_SD_CARD_NIOS_timer;

	component DE2_115_SD_CARD_NIOS_tri_state_bridge_flash_bridge_0 is
		port (
			clk                                   : in    std_logic                     := 'X';             -- clk
			reset                                 : in    std_logic                     := 'X';             -- reset
			request                               : in    std_logic                     := 'X';             -- request
			grant                                 : out   std_logic;                                        -- grant
			tcs_address_to_the_cfi_flash          : in    std_logic_vector(22 downto 0) := (others => 'X'); -- address_to_the_cfi_flash_out
			tcs_tri_state_bridge_flash_data       : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_flash_data_out
			tcs_tri_state_bridge_flash_data_outen : in    std_logic                     := 'X';             -- tri_state_bridge_flash_data_outen
			tcs_tri_state_bridge_flash_data_in    : out   std_logic_vector(7 downto 0);                     -- tri_state_bridge_flash_data_in
			tcs_write_n_to_the_cfi_flash          : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_to_the_cfi_flash_out
			tcs_select_n_to_the_cfi_flash         : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- select_n_to_the_cfi_flash_out
			tcs_read_n_to_the_cfi_flash           : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- read_n_to_the_cfi_flash_out
			address_to_the_cfi_flash              : out   std_logic_vector(22 downto 0);                    -- address_to_the_cfi_flash
			tri_state_bridge_flash_data           : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_flash_data
			write_n_to_the_cfi_flash              : out   std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash
			select_n_to_the_cfi_flash             : out   std_logic_vector(0 downto 0);                     -- select_n_to_the_cfi_flash
			read_n_to_the_cfi_flash               : out   std_logic_vector(0 downto 0)                      -- read_n_to_the_cfi_flash
		);
	end component DE2_115_SD_CARD_NIOS_tri_state_bridge_flash_bridge_0;

	component DE2_115_SD_CARD_NIOS_tri_state_flash_bridge_pinSharer_0 is
		port (
			clk_clk                           : in  std_logic                     := 'X';             -- clk
			reset_reset                       : in  std_logic                     := 'X';             -- reset
			request                           : out std_logic;                                        -- request
			grant                             : in  std_logic                     := 'X';             -- grant
			address_to_the_cfi_flash          : out std_logic_vector(22 downto 0);                    -- address_to_the_cfi_flash_out
			read_n_to_the_cfi_flash           : out std_logic_vector(0 downto 0);                     -- read_n_to_the_cfi_flash_out
			write_n_to_the_cfi_flash          : out std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash_out
			tri_state_bridge_flash_data       : out std_logic_vector(7 downto 0);                     -- tri_state_bridge_flash_data_out
			tri_state_bridge_flash_data_in    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_flash_data_in
			tri_state_bridge_flash_data_outen : out std_logic;                                        -- tri_state_bridge_flash_data_outen
			select_n_to_the_cfi_flash         : out std_logic_vector(0 downto 0);                     -- select_n_to_the_cfi_flash_out
			tcs0_request                      : in  std_logic                     := 'X';             -- request
			tcs0_grant                        : out std_logic;                                        -- grant
			tcs0_address_out                  : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address_out
			tcs0_read_n_out                   : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- read_n_out
			tcs0_write_n_out                  : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs0_data_out                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_out
			tcs0_data_in                      : out std_logic_vector(7 downto 0);                     -- data_in
			tcs0_data_outen                   : in  std_logic                     := 'X';             -- data_outen
			tcs0_chipselect_n_out             : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- chipselect_n_out
		);
	end component DE2_115_SD_CARD_NIOS_tri_state_flash_bridge_pinSharer_0;

	component DE2_115_SD_CARD_NIOS_video_character_buffer_with_dma_0 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			ctrl_address         : in  std_logic                     := 'X';             -- address
			ctrl_byteenable      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ctrl_chipselect      : in  std_logic                     := 'X';             -- chipselect
			ctrl_read            : in  std_logic                     := 'X';             -- read
			ctrl_write           : in  std_logic                     := 'X';             -- write
			ctrl_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ctrl_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			buf_byteenable       : in  std_logic                     := 'X';             -- byteenable
			buf_chipselect       : in  std_logic                     := 'X';             -- chipselect
			buf_read             : in  std_logic                     := 'X';             -- read
			buf_write            : in  std_logic                     := 'X';             -- write
			buf_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			buf_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			buf_waitrequest      : out std_logic;                                        -- waitrequest
			buf_address          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component DE2_115_SD_CARD_NIOS_video_character_buffer_with_dma_0;

	component DE2_115_SD_CARD_NIOS_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			lcd_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component DE2_115_SD_CARD_NIOS_video_pll_0;

	component DE2_115_SD_CARD_NIOS_video_vga_controller_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component DE2_115_SD_CARD_NIOS_video_vga_controller_0;

	component DE2_115_SD_CARD_NIOS_weight_index is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(12 downto 0)                     -- export
		);
	end component DE2_115_SD_CARD_NIOS_weight_index;

	component DE2_115_SD_CARD_NIOS_mm_interconnect_0 is
		port (
			altpll_c0_clk                                                          : in  std_logic                     := 'X';             -- clk
			clk_50_clk_clk                                                         : in  std_logic                     := 'X';             -- clk
			video_pll_0_vga_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			altpll_inclk_interface_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			cpu_reset_reset_bridge_in_reset_reset                                  : in  std_logic                     := 'X';             -- reset
			onchip_memory2_reset1_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			video_character_buffer_with_dma_0_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                                : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                            : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                                   : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                               : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid                                          : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                                                  : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                            : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                                         : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                                     : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                                            : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                                        : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                                   : out std_logic;                                        -- readdatavalid
			activations_index_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			activations_index_s1_write                                             : out std_logic;                                        -- write
			activations_index_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			activations_index_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			activations_index_s1_chipselect                                        : out std_logic;                                        -- chipselect
			altpll_pll_slave_address                                               : out std_logic_vector(1 downto 0);                     -- address
			altpll_pll_slave_write                                                 : out std_logic;                                        -- write
			altpll_pll_slave_read                                                  : out std_logic;                                        -- read
			altpll_pll_slave_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_pll_slave_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			cfi_flash_uas_address                                                  : out std_logic_vector(22 downto 0);                    -- address
			cfi_flash_uas_write                                                    : out std_logic;                                        -- write
			cfi_flash_uas_read                                                     : out std_logic;                                        -- read
			cfi_flash_uas_readdata                                                 : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			cfi_flash_uas_writedata                                                : out std_logic_vector(7 downto 0);                     -- writedata
			cfi_flash_uas_burstcount                                               : out std_logic_vector(0 downto 0);                     -- burstcount
			cfi_flash_uas_byteenable                                               : out std_logic_vector(0 downto 0);                     -- byteenable
			cfi_flash_uas_readdatavalid                                            : in  std_logic                     := 'X';             -- readdatavalid
			cfi_flash_uas_waitrequest                                              : in  std_logic                     := 'X';             -- waitrequest
			cfi_flash_uas_lock                                                     : out std_logic;                                        -- lock
			cfi_flash_uas_debugaccess                                              : out std_logic;                                        -- debugaccess
			clock_crossing_io_s0_address                                           : out std_logic_vector(8 downto 0);                     -- address
			clock_crossing_io_s0_write                                             : out std_logic;                                        -- write
			clock_crossing_io_s0_read                                              : out std_logic;                                        -- read
			clock_crossing_io_s0_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			clock_crossing_io_s0_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			clock_crossing_io_s0_burstcount                                        : out std_logic_vector(0 downto 0);                     -- burstcount
			clock_crossing_io_s0_byteenable                                        : out std_logic_vector(3 downto 0);                     -- byteenable
			clock_crossing_io_s0_readdatavalid                                     : in  std_logic                     := 'X';             -- readdatavalid
			clock_crossing_io_s0_waitrequest                                       : in  std_logic                     := 'X';             -- waitrequest
			clock_crossing_io_s0_debugaccess                                       : out std_logic;                                        -- debugaccess
			cpu_debug_mem_slave_address                                            : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                              : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                               : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                                         : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                                        : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                                        : out std_logic;                                        -- debugaccess
			floatdata_output_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			floatdata_output_s1_write                                              : out std_logic;                                        -- write
			floatdata_output_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			floatdata_output_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			floatdata_output_s1_chipselect                                         : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                                    : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                                      : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                                       : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                                : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                                 : out std_logic;                                        -- chipselect
			key_s1_address                                                         : out std_logic_vector(1 downto 0);                     -- address
			key_s1_write                                                           : out std_logic;                                        -- write
			key_s1_readdata                                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_s1_writedata                                                       : out std_logic_vector(31 downto 0);                    -- writedata
			key_s1_chipselect                                                      : out std_logic;                                        -- chipselect
			ledg_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			ledg_s1_write                                                          : out std_logic;                                        -- write
			ledg_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ledg_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			ledg_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			ledr_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			ledr_s1_write                                                          : out std_logic;                                        -- write
			ledr_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ledr_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			ledr_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			onchip_memory2_s1_address                                              : out std_logic_vector(15 downto 0);                    -- address
			onchip_memory2_s1_write                                                : out std_logic;                                        -- write
			onchip_memory2_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_s1_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_s1_byteenable                                           : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_s1_chipselect                                           : out std_logic;                                        -- chipselect
			onchip_memory2_s1_clken                                                : out std_logic;                                        -- clken
			pixel_index_s1_address                                                 : out std_logic_vector(1 downto 0);                     -- address
			pixel_index_s1_write                                                   : out std_logic;                                        -- write
			pixel_index_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pixel_index_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			pixel_index_s1_chipselect                                              : out std_logic;                                        -- chipselect
			results_input_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			results_input_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sw_s1_address                                                          : out std_logic_vector(1 downto 0);                     -- address
			sw_s1_write                                                            : out std_logic;                                        -- write
			sw_s1_readdata                                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sw_s1_writedata                                                        : out std_logic_vector(31 downto 0);                    -- writedata
			sw_s1_chipselect                                                       : out std_logic;                                        -- chipselect
			sync_data_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			sync_data_s1_write                                                     : out std_logic;                                        -- write
			sync_data_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sync_data_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			sync_data_s1_chipselect                                                : out std_logic;                                        -- chipselect
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     : out std_logic_vector(12 downto 0);                    -- address
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       : out std_logic;                                        -- write
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        : out std_logic;                                        -- read
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  : out std_logic_vector(0 downto 0);                     -- byteenable
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  : out std_logic;                                        -- chipselect
			video_character_buffer_with_dma_0_avalon_char_control_slave_address    : out std_logic_vector(0 downto 0);                     -- address
			video_character_buffer_with_dma_0_avalon_char_control_slave_write      : out std_logic;                                        -- write
			video_character_buffer_with_dma_0_avalon_char_control_slave_read       : out std_logic;                                        -- read
			video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable : out std_logic_vector(3 downto 0);                     -- byteenable
			video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect : out std_logic;                                        -- chipselect
			weight_index_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			weight_index_s1_write                                                  : out std_logic;                                        -- write
			weight_index_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			weight_index_s1_writedata                                              : out std_logic_vector(31 downto 0);                    -- writedata
			weight_index_s1_chipselect                                             : out std_logic                                         -- chipselect
		);
	end component DE2_115_SD_CARD_NIOS_mm_interconnect_0;

	component DE2_115_SD_CARD_NIOS_mm_interconnect_1 is
		port (
			altpll_c0_clk                                          : in  std_logic                     := 'X';             -- clk
			altpll_c2_clk                                          : in  std_logic                     := 'X';             -- clk
			clock_crossing_io_m0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sd_clk_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			clock_crossing_io_m0_address                           : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			clock_crossing_io_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			clock_crossing_io_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			clock_crossing_io_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock_crossing_io_m0_read                              : in  std_logic                     := 'X';             -- read
			clock_crossing_io_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			clock_crossing_io_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			clock_crossing_io_m0_write                             : in  std_logic                     := 'X';             -- write
			clock_crossing_io_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_crossing_io_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			sd_clk_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			sd_clk_s1_write                                        : out std_logic;                                        -- write
			sd_clk_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sd_clk_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			sd_clk_s1_chipselect                                   : out std_logic;                                        -- chipselect
			sd_cmd_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			sd_cmd_s1_write                                        : out std_logic;                                        -- write
			sd_cmd_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sd_cmd_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			sd_cmd_s1_chipselect                                   : out std_logic;                                        -- chipselect
			sd_dat_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			sd_dat_s1_write                                        : out std_logic;                                        -- write
			sd_dat_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sd_dat_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			sd_dat_s1_chipselect                                   : out std_logic;                                        -- chipselect
			sd_wp_n_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			sd_wp_n_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                                       : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                                         : out std_logic;                                        -- write
			timer_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                                    : out std_logic                                         -- chipselect
		);
	end component DE2_115_SD_CARD_NIOS_mm_interconnect_1;

	component DE2_115_SD_CARD_NIOS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DE2_115_SD_CARD_NIOS_irq_mapper;

	component de2_115_sd_card_nios_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de2_115_sd_card_nios_rst_controller;

	component de2_115_sd_card_nios_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de2_115_sd_card_nios_rst_controller_001;

	component de2_115_sd_card_nios_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de2_115_sd_card_nios_rst_controller_002;

	component de2_115_sd_card_nios_rst_controller_004 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de2_115_sd_card_nios_rst_controller_004;

	signal video_character_buffer_with_dma_0_avalon_char_source_valid                               : std_logic;                     -- video_character_buffer_with_dma_0:stream_valid -> video_vga_controller_0:valid
	signal video_character_buffer_with_dma_0_avalon_char_source_data                                : std_logic_vector(29 downto 0); -- video_character_buffer_with_dma_0:stream_data -> video_vga_controller_0:data
	signal video_character_buffer_with_dma_0_avalon_char_source_ready                               : std_logic;                     -- video_vga_controller_0:ready -> video_character_buffer_with_dma_0:stream_ready
	signal video_character_buffer_with_dma_0_avalon_char_source_startofpacket                       : std_logic;                     -- video_character_buffer_with_dma_0:stream_startofpacket -> video_vga_controller_0:startofpacket
	signal video_character_buffer_with_dma_0_avalon_char_source_endofpacket                         : std_logic;                     -- video_character_buffer_with_dma_0:stream_endofpacket -> video_vga_controller_0:endofpacket
	signal altpll_c0_clk                                                                            : std_logic;                     -- altpll:c0 -> [c0_out_clk_clk, activations_index:clk, cfi_flash:clk_clk, clock_crossing_io:s0_clk, cpu:clk, floatdata_output:clk, irq_mapper:clk, jtag_uart:clk, key:clk, ledg:clk, ledr:clk, mm_interconnect_0:altpll_c0_clk, mm_interconnect_1:altpll_c0_clk, onchip_memory2:clk, pixel_index:clk, results_input:clk, rst_controller:clk, rst_controller_002:clk, sd_clk:clk, sd_cmd:clk, sd_dat:clk, sd_wp_n:clk, sw:clk, sync_data:clk, timer:clk, tri_state_bridge_flash_bridge_0:clk, tri_state_flash_bridge_pinSharer_0:clk_clk, weight_index:clk]
	signal altpll_c2_clk                                                                            : std_logic;                     -- altpll:c2 -> [c2_out_clk_clk, clock_crossing_io:m0_clk, mm_interconnect_1:altpll_c2_clk, rst_controller_003:clk]
	signal video_pll_0_vga_clk_clk                                                                  : std_logic;                     -- video_pll_0:vga_clk_clk -> [mm_interconnect_0:video_pll_0_vga_clk_clk, rst_controller_004:clk, video_character_buffer_with_dma_0:clk, video_vga_controller_0:clk]
	signal tri_state_flash_bridge_pinsharer_0_tcm_request                                           : std_logic;                     -- tri_state_flash_bridge_pinSharer_0:request -> tri_state_bridge_flash_bridge_0:request
	signal tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out                       : std_logic_vector(0 downto 0);  -- tri_state_flash_bridge_pinSharer_0:read_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_read_n_to_the_cfi_flash
	signal tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out                      : std_logic_vector(22 downto 0); -- tri_state_flash_bridge_pinSharer_0:address_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_address_to_the_cfi_flash
	signal tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen                 : std_logic;                     -- tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data_outen -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_outen
	signal tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out                      : std_logic_vector(0 downto 0);  -- tri_state_flash_bridge_pinSharer_0:write_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_write_n_to_the_cfi_flash
	signal tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in                    : std_logic_vector(7 downto 0);  -- tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_in -> tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data_in
	signal tri_state_flash_bridge_pinsharer_0_tcm_grant                                             : std_logic;                     -- tri_state_bridge_flash_bridge_0:grant -> tri_state_flash_bridge_pinSharer_0:grant
	signal tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out                   : std_logic_vector(7 downto 0);  -- tri_state_flash_bridge_pinSharer_0:tri_state_bridge_flash_data -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data
	signal tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out                     : std_logic_vector(0 downto 0);  -- tri_state_flash_bridge_pinSharer_0:select_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_select_n_to_the_cfi_flash
	signal cfi_flash_tcm_data_outen                                                                 : std_logic;                     -- cfi_flash:tcm_data_outen -> tri_state_flash_bridge_pinSharer_0:tcs0_data_outen
	signal cfi_flash_tcm_request                                                                    : std_logic;                     -- cfi_flash:tcm_request -> tri_state_flash_bridge_pinSharer_0:tcs0_request
	signal cfi_flash_tcm_write_n_out                                                                : std_logic;                     -- cfi_flash:tcm_write_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_write_n_out
	signal cfi_flash_tcm_read_n_out                                                                 : std_logic;                     -- cfi_flash:tcm_read_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_read_n_out
	signal cfi_flash_tcm_grant                                                                      : std_logic;                     -- tri_state_flash_bridge_pinSharer_0:tcs0_grant -> cfi_flash:tcm_grant
	signal cfi_flash_tcm_chipselect_n_out                                                           : std_logic;                     -- cfi_flash:tcm_chipselect_n_out -> tri_state_flash_bridge_pinSharer_0:tcs0_chipselect_n_out
	signal cfi_flash_tcm_address_out                                                                : std_logic_vector(22 downto 0); -- cfi_flash:tcm_address_out -> tri_state_flash_bridge_pinSharer_0:tcs0_address_out
	signal cfi_flash_tcm_data_out                                                                   : std_logic_vector(7 downto 0);  -- cfi_flash:tcm_data_out -> tri_state_flash_bridge_pinSharer_0:tcs0_data_out
	signal cfi_flash_tcm_data_in                                                                    : std_logic_vector(7 downto 0);  -- tri_state_flash_bridge_pinSharer_0:tcs0_data_in -> cfi_flash:tcm_data_in
	signal cpu_data_master_readdata                                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                                              : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                                              : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                                  : std_logic_vector(25 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                               : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                                     : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                                            : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                                                    : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                                : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                                       : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                                           : std_logic_vector(25 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                                              : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                                                     : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    : std_logic_vector(7 downto 0);  -- video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest : std_logic;                     -- video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     : std_logic_vector(12 downto 0); -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   : std_logic_vector(7 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   : std_logic_vector(31 downto 0); -- video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read       : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write      : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect                                 : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                                   : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest                                : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                                    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                                       : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                                      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                                           : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                                        : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                                        : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                                            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                               : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                                              : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_pll_slave_readdata                                              : std_logic_vector(31 downto 0); -- altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	signal mm_interconnect_0_altpll_pll_slave_address                                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	signal mm_interconnect_0_altpll_pll_slave_read                                                  : std_logic;                     -- mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	signal mm_interconnect_0_altpll_pll_slave_write                                                 : std_logic;                     -- mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	signal mm_interconnect_0_altpll_pll_slave_writedata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	signal mm_interconnect_0_clock_crossing_io_s0_readdata                                          : std_logic_vector(31 downto 0); -- clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	signal mm_interconnect_0_clock_crossing_io_s0_waitrequest                                       : std_logic;                     -- clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	signal mm_interconnect_0_clock_crossing_io_s0_debugaccess                                       : std_logic;                     -- mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	signal mm_interconnect_0_clock_crossing_io_s0_address                                           : std_logic_vector(8 downto 0);  -- mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	signal mm_interconnect_0_clock_crossing_io_s0_read                                              : std_logic;                     -- mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	signal mm_interconnect_0_clock_crossing_io_s0_byteenable                                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	signal mm_interconnect_0_clock_crossing_io_s0_readdatavalid                                     : std_logic;                     -- clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	signal mm_interconnect_0_clock_crossing_io_s0_write                                             : std_logic;                     -- mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	signal mm_interconnect_0_clock_crossing_io_s0_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	signal mm_interconnect_0_clock_crossing_io_s0_burstcount                                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	signal mm_interconnect_0_onchip_memory2_s1_chipselect                                           : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	signal mm_interconnect_0_onchip_memory2_s1_readdata                                             : std_logic_vector(31 downto 0); -- onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	signal mm_interconnect_0_onchip_memory2_s1_address                                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	signal mm_interconnect_0_onchip_memory2_s1_byteenable                                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	signal mm_interconnect_0_onchip_memory2_s1_write                                                : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	signal mm_interconnect_0_onchip_memory2_s1_writedata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	signal mm_interconnect_0_onchip_memory2_s1_clken                                                : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	signal mm_interconnect_0_ledr_s1_chipselect                                                     : std_logic;                     -- mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	signal mm_interconnect_0_ledr_s1_readdata                                                       : std_logic_vector(31 downto 0); -- ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	signal mm_interconnect_0_ledr_s1_address                                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ledr_s1_address -> ledr:address
	signal mm_interconnect_0_ledr_s1_write                                                          : std_logic;                     -- mm_interconnect_0:ledr_s1_write -> mm_interconnect_0_ledr_s1_write:in
	signal mm_interconnect_0_ledr_s1_writedata                                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	signal mm_interconnect_0_ledg_s1_chipselect                                                     : std_logic;                     -- mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	signal mm_interconnect_0_ledg_s1_readdata                                                       : std_logic_vector(31 downto 0); -- ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	signal mm_interconnect_0_ledg_s1_address                                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ledg_s1_address -> ledg:address
	signal mm_interconnect_0_ledg_s1_write                                                          : std_logic;                     -- mm_interconnect_0:ledg_s1_write -> mm_interconnect_0_ledg_s1_write:in
	signal mm_interconnect_0_ledg_s1_writedata                                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	signal mm_interconnect_0_sw_s1_chipselect                                                       : std_logic;                     -- mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	signal mm_interconnect_0_sw_s1_readdata                                                         : std_logic_vector(31 downto 0); -- sw:readdata -> mm_interconnect_0:sw_s1_readdata
	signal mm_interconnect_0_sw_s1_address                                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sw_s1_address -> sw:address
	signal mm_interconnect_0_sw_s1_write                                                            : std_logic;                     -- mm_interconnect_0:sw_s1_write -> mm_interconnect_0_sw_s1_write:in
	signal mm_interconnect_0_sw_s1_writedata                                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sw_s1_writedata -> sw:writedata
	signal mm_interconnect_0_key_s1_chipselect                                                      : std_logic;                     -- mm_interconnect_0:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_0_key_s1_readdata                                                        : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_key_s1_write                                                           : std_logic;                     -- mm_interconnect_0:key_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_writedata                                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_s1_writedata -> key:writedata
	signal mm_interconnect_0_floatdata_output_s1_chipselect                                         : std_logic;                     -- mm_interconnect_0:floatdata_output_s1_chipselect -> floatdata_output:chipselect
	signal mm_interconnect_0_floatdata_output_s1_readdata                                           : std_logic_vector(31 downto 0); -- floatdata_output:readdata -> mm_interconnect_0:floatdata_output_s1_readdata
	signal mm_interconnect_0_floatdata_output_s1_address                                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:floatdata_output_s1_address -> floatdata_output:address
	signal mm_interconnect_0_floatdata_output_s1_write                                              : std_logic;                     -- mm_interconnect_0:floatdata_output_s1_write -> mm_interconnect_0_floatdata_output_s1_write:in
	signal mm_interconnect_0_floatdata_output_s1_writedata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:floatdata_output_s1_writedata -> floatdata_output:writedata
	signal mm_interconnect_0_sync_data_s1_chipselect                                                : std_logic;                     -- mm_interconnect_0:sync_data_s1_chipselect -> sync_data:chipselect
	signal mm_interconnect_0_sync_data_s1_readdata                                                  : std_logic_vector(31 downto 0); -- sync_data:readdata -> mm_interconnect_0:sync_data_s1_readdata
	signal mm_interconnect_0_sync_data_s1_address                                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sync_data_s1_address -> sync_data:address
	signal mm_interconnect_0_sync_data_s1_write                                                     : std_logic;                     -- mm_interconnect_0:sync_data_s1_write -> mm_interconnect_0_sync_data_s1_write:in
	signal mm_interconnect_0_sync_data_s1_writedata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:sync_data_s1_writedata -> sync_data:writedata
	signal mm_interconnect_0_pixel_index_s1_chipselect                                              : std_logic;                     -- mm_interconnect_0:pixel_index_s1_chipselect -> pixel_index:chipselect
	signal mm_interconnect_0_pixel_index_s1_readdata                                                : std_logic_vector(31 downto 0); -- pixel_index:readdata -> mm_interconnect_0:pixel_index_s1_readdata
	signal mm_interconnect_0_pixel_index_s1_address                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pixel_index_s1_address -> pixel_index:address
	signal mm_interconnect_0_pixel_index_s1_write                                                   : std_logic;                     -- mm_interconnect_0:pixel_index_s1_write -> mm_interconnect_0_pixel_index_s1_write:in
	signal mm_interconnect_0_pixel_index_s1_writedata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:pixel_index_s1_writedata -> pixel_index:writedata
	signal mm_interconnect_0_weight_index_s1_chipselect                                             : std_logic;                     -- mm_interconnect_0:weight_index_s1_chipselect -> weight_index:chipselect
	signal mm_interconnect_0_weight_index_s1_readdata                                               : std_logic_vector(31 downto 0); -- weight_index:readdata -> mm_interconnect_0:weight_index_s1_readdata
	signal mm_interconnect_0_weight_index_s1_address                                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:weight_index_s1_address -> weight_index:address
	signal mm_interconnect_0_weight_index_s1_write                                                  : std_logic;                     -- mm_interconnect_0:weight_index_s1_write -> mm_interconnect_0_weight_index_s1_write:in
	signal mm_interconnect_0_weight_index_s1_writedata                                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:weight_index_s1_writedata -> weight_index:writedata
	signal mm_interconnect_0_results_input_s1_readdata                                              : std_logic_vector(31 downto 0); -- results_input:readdata -> mm_interconnect_0:results_input_s1_readdata
	signal mm_interconnect_0_results_input_s1_address                                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:results_input_s1_address -> results_input:address
	signal mm_interconnect_0_activations_index_s1_chipselect                                        : std_logic;                     -- mm_interconnect_0:activations_index_s1_chipselect -> activations_index:chipselect
	signal mm_interconnect_0_activations_index_s1_readdata                                          : std_logic_vector(31 downto 0); -- activations_index:readdata -> mm_interconnect_0:activations_index_s1_readdata
	signal mm_interconnect_0_activations_index_s1_address                                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:activations_index_s1_address -> activations_index:address
	signal mm_interconnect_0_activations_index_s1_write                                             : std_logic;                     -- mm_interconnect_0:activations_index_s1_write -> mm_interconnect_0_activations_index_s1_write:in
	signal mm_interconnect_0_activations_index_s1_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:activations_index_s1_writedata -> activations_index:writedata
	signal mm_interconnect_0_cfi_flash_uas_readdata                                                 : std_logic_vector(7 downto 0);  -- cfi_flash:uas_readdata -> mm_interconnect_0:cfi_flash_uas_readdata
	signal mm_interconnect_0_cfi_flash_uas_waitrequest                                              : std_logic;                     -- cfi_flash:uas_waitrequest -> mm_interconnect_0:cfi_flash_uas_waitrequest
	signal mm_interconnect_0_cfi_flash_uas_debugaccess                                              : std_logic;                     -- mm_interconnect_0:cfi_flash_uas_debugaccess -> cfi_flash:uas_debugaccess
	signal mm_interconnect_0_cfi_flash_uas_address                                                  : std_logic_vector(22 downto 0); -- mm_interconnect_0:cfi_flash_uas_address -> cfi_flash:uas_address
	signal mm_interconnect_0_cfi_flash_uas_read                                                     : std_logic;                     -- mm_interconnect_0:cfi_flash_uas_read -> cfi_flash:uas_read
	signal mm_interconnect_0_cfi_flash_uas_byteenable                                               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:cfi_flash_uas_byteenable -> cfi_flash:uas_byteenable
	signal mm_interconnect_0_cfi_flash_uas_readdatavalid                                            : std_logic;                     -- cfi_flash:uas_readdatavalid -> mm_interconnect_0:cfi_flash_uas_readdatavalid
	signal mm_interconnect_0_cfi_flash_uas_lock                                                     : std_logic;                     -- mm_interconnect_0:cfi_flash_uas_lock -> cfi_flash:uas_lock
	signal mm_interconnect_0_cfi_flash_uas_write                                                    : std_logic;                     -- mm_interconnect_0:cfi_flash_uas_write -> cfi_flash:uas_write
	signal mm_interconnect_0_cfi_flash_uas_writedata                                                : std_logic_vector(7 downto 0);  -- mm_interconnect_0:cfi_flash_uas_writedata -> cfi_flash:uas_writedata
	signal mm_interconnect_0_cfi_flash_uas_burstcount                                               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:cfi_flash_uas_burstcount -> cfi_flash:uas_burstcount
	signal clock_crossing_io_m0_waitrequest                                                         : std_logic;                     -- mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	signal clock_crossing_io_m0_readdata                                                            : std_logic_vector(31 downto 0); -- mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	signal clock_crossing_io_m0_debugaccess                                                         : std_logic;                     -- clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	signal clock_crossing_io_m0_address                                                             : std_logic_vector(8 downto 0);  -- clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	signal clock_crossing_io_m0_read                                                                : std_logic;                     -- clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	signal clock_crossing_io_m0_byteenable                                                          : std_logic_vector(3 downto 0);  -- clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	signal clock_crossing_io_m0_readdatavalid                                                       : std_logic;                     -- mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	signal clock_crossing_io_m0_writedata                                                           : std_logic_vector(31 downto 0); -- clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	signal clock_crossing_io_m0_write                                                               : std_logic;                     -- clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	signal clock_crossing_io_m0_burstcount                                                          : std_logic_vector(0 downto 0);  -- clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	signal mm_interconnect_1_sd_clk_s1_chipselect                                                   : std_logic;                     -- mm_interconnect_1:sd_clk_s1_chipselect -> sd_clk:chipselect
	signal mm_interconnect_1_sd_clk_s1_readdata                                                     : std_logic_vector(31 downto 0); -- sd_clk:readdata -> mm_interconnect_1:sd_clk_s1_readdata
	signal mm_interconnect_1_sd_clk_s1_address                                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sd_clk_s1_address -> sd_clk:address
	signal mm_interconnect_1_sd_clk_s1_write                                                        : std_logic;                     -- mm_interconnect_1:sd_clk_s1_write -> mm_interconnect_1_sd_clk_s1_write:in
	signal mm_interconnect_1_sd_clk_s1_writedata                                                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:sd_clk_s1_writedata -> sd_clk:writedata
	signal mm_interconnect_1_sd_cmd_s1_chipselect                                                   : std_logic;                     -- mm_interconnect_1:sd_cmd_s1_chipselect -> sd_cmd:chipselect
	signal mm_interconnect_1_sd_cmd_s1_readdata                                                     : std_logic_vector(31 downto 0); -- sd_cmd:readdata -> mm_interconnect_1:sd_cmd_s1_readdata
	signal mm_interconnect_1_sd_cmd_s1_address                                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sd_cmd_s1_address -> sd_cmd:address
	signal mm_interconnect_1_sd_cmd_s1_write                                                        : std_logic;                     -- mm_interconnect_1:sd_cmd_s1_write -> mm_interconnect_1_sd_cmd_s1_write:in
	signal mm_interconnect_1_sd_cmd_s1_writedata                                                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:sd_cmd_s1_writedata -> sd_cmd:writedata
	signal mm_interconnect_1_sd_dat_s1_chipselect                                                   : std_logic;                     -- mm_interconnect_1:sd_dat_s1_chipselect -> sd_dat:chipselect
	signal mm_interconnect_1_sd_dat_s1_readdata                                                     : std_logic_vector(31 downto 0); -- sd_dat:readdata -> mm_interconnect_1:sd_dat_s1_readdata
	signal mm_interconnect_1_sd_dat_s1_address                                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sd_dat_s1_address -> sd_dat:address
	signal mm_interconnect_1_sd_dat_s1_write                                                        : std_logic;                     -- mm_interconnect_1:sd_dat_s1_write -> mm_interconnect_1_sd_dat_s1_write:in
	signal mm_interconnect_1_sd_dat_s1_writedata                                                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:sd_dat_s1_writedata -> sd_dat:writedata
	signal mm_interconnect_1_sd_wp_n_s1_readdata                                                    : std_logic_vector(31 downto 0); -- sd_wp_n:readdata -> mm_interconnect_1:sd_wp_n_s1_readdata
	signal mm_interconnect_1_sd_wp_n_s1_address                                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sd_wp_n_s1_address -> sd_wp_n:address
	signal mm_interconnect_1_timer_s1_chipselect                                                    : std_logic;                     -- mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_1_timer_s1_readdata                                                      : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_1:timer_s1_readdata
	signal mm_interconnect_1_timer_s1_address                                                       : std_logic_vector(2 downto 0);  -- mm_interconnect_1:timer_s1_address -> timer:address
	signal mm_interconnect_1_timer_s1_write                                                         : std_logic;                     -- mm_interconnect_1:timer_s1_write -> mm_interconnect_1_timer_s1_write:in
	signal mm_interconnect_1_timer_s1_writedata                                                     : std_logic_vector(15 downto 0); -- mm_interconnect_1:timer_s1_writedata -> timer:writedata
	signal irq_mapper_receiver0_irq                                                                 : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                 : std_logic;                     -- timer:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                                           : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:onchip_memory2_reset1_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                                       : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                                       : std_logic;                     -- rst_controller_001:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal cpu_debug_reset_request_reset                                                            : std_logic;                     -- cpu:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	signal rst_controller_002_reset_out_reset                                                       : std_logic;                     -- rst_controller_002:reset_out -> [cfi_flash:reset_reset, clock_crossing_io:s0_reset, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sd_clk_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in, rst_translator_001:in_reset, tri_state_bridge_flash_bridge_0:reset, tri_state_flash_bridge_pinSharer_0:reset_reset]
	signal rst_controller_002_reset_out_reset_req                                                   : std_logic;                     -- rst_controller_002:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_003_reset_out_reset                                                       : std_logic;                     -- rst_controller_003:reset_out -> [clock_crossing_io:m0_reset, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset]
	signal rst_controller_004_reset_out_reset                                                       : std_logic;                     -- rst_controller_004:reset_out -> [mm_interconnect_0:video_character_buffer_with_dma_0_reset_reset_bridge_in_reset_reset, video_character_buffer_with_dma_0:reset, video_vga_controller_0:reset]
	signal video_pll_0_reset_source_reset                                                           : std_logic;                     -- video_pll_0:reset_source_reset -> rst_controller_004:reset_in0
	signal rst_controller_005_reset_out_reset                                                       : std_logic;                     -- rst_controller_005:reset_out -> video_pll_0:ref_reset_reset
	signal reset_reset_n_ports_inv                                                                  : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_005:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv                             : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_ledr_s1_write_ports_inv                                                : std_logic;                     -- mm_interconnect_0_ledr_s1_write:inv -> ledr:write_n
	signal mm_interconnect_0_ledg_s1_write_ports_inv                                                : std_logic;                     -- mm_interconnect_0_ledg_s1_write:inv -> ledg:write_n
	signal mm_interconnect_0_sw_s1_write_ports_inv                                                  : std_logic;                     -- mm_interconnect_0_sw_s1_write:inv -> sw:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                                                 : std_logic;                     -- mm_interconnect_0_key_s1_write:inv -> key:write_n
	signal mm_interconnect_0_floatdata_output_s1_write_ports_inv                                    : std_logic;                     -- mm_interconnect_0_floatdata_output_s1_write:inv -> floatdata_output:write_n
	signal mm_interconnect_0_sync_data_s1_write_ports_inv                                           : std_logic;                     -- mm_interconnect_0_sync_data_s1_write:inv -> sync_data:write_n
	signal mm_interconnect_0_pixel_index_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_0_pixel_index_s1_write:inv -> pixel_index:write_n
	signal mm_interconnect_0_weight_index_s1_write_ports_inv                                        : std_logic;                     -- mm_interconnect_0_weight_index_s1_write:inv -> weight_index:write_n
	signal mm_interconnect_0_activations_index_s1_write_ports_inv                                   : std_logic;                     -- mm_interconnect_0_activations_index_s1_write:inv -> activations_index:write_n
	signal mm_interconnect_1_sd_clk_s1_write_ports_inv                                              : std_logic;                     -- mm_interconnect_1_sd_clk_s1_write:inv -> sd_clk:write_n
	signal mm_interconnect_1_sd_cmd_s1_write_ports_inv                                              : std_logic;                     -- mm_interconnect_1_sd_cmd_s1_write:inv -> sd_cmd:write_n
	signal mm_interconnect_1_sd_dat_s1_write_ports_inv                                              : std_logic;                     -- mm_interconnect_1_sd_dat_s1_write:inv -> sd_dat:write_n
	signal mm_interconnect_1_timer_s1_write_ports_inv                                               : std_logic;                     -- mm_interconnect_1_timer_s1_write:inv -> timer:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [activations_index:reset_n, floatdata_output:reset_n, key:reset_n, ledg:reset_n, ledr:reset_n, pixel_index:reset_n, results_input:reset_n, sw:reset_n, sync_data:reset_n, weight_index:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                                             : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n, sd_clk:reset_n, sd_cmd:reset_n, sd_dat:reset_n, sd_wp_n:reset_n, timer:reset_n]

begin

	activations_index : component DE2_115_SD_CARD_NIOS_activations_index
		port map (
			clk        => altpll_c0_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,               --               reset.reset_n
			address    => mm_interconnect_0_activations_index_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_activations_index_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_activations_index_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_activations_index_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_activations_index_s1_readdata,        --                    .readdata
			out_port   => activations_index_external_connection_export            -- external_connection.export
		);

	altpll : component DE2_115_SD_CARD_NIOS_altpll
		port map (
			clk                => clk_50_clk_in_clk,                            --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,           -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_pll_slave_writedata, --                      .writedata
			c0                 => altpll_c0_clk,                                --                    c0.clk
			c1                 => altpll_c1_clk,                                --                    c1.clk
			c2                 => altpll_c2_clk,                                --                    c2.clk
			c3                 => altpll_c3_clk,                                --                    c3.clk
			areset             => altpll_areset_conduit_export,                 --        areset_conduit.export
			locked             => altpll_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                         --           (terminated)
			scandataout        => open,                                         --           (terminated)
			phasecounterselect => "0000",                                       --           (terminated)
			phaseupdown        => '0',                                          --           (terminated)
			phasestep          => '0',                                          --           (terminated)
			scanclk            => '0',                                          --           (terminated)
			scanclkena         => '0',                                          --           (terminated)
			scandata           => '0',                                          --           (terminated)
			configupdate       => '0',                                          --           (terminated)
			phasedone          => open                                          --           (terminated)
		);

	cfi_flash : component DE2_115_SD_CARD_NIOS_cfi_flash
		generic map (
			TCM_ADDRESS_W                  => 23,
			TCM_DATA_W                     => 8,
			TCM_BYTEENABLE_W               => 1,
			TCM_READ_WAIT                  => 0,
			TCM_WRITE_WAIT                 => 0,
			TCM_SETUP_WAIT                 => 0,
			TCM_DATA_HOLD                  => 0,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 1,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => altpll_c0_clk,                                 --   clk.clk
			reset_reset          => rst_controller_002_reset_out_reset,            -- reset.reset
			uas_address          => mm_interconnect_0_cfi_flash_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_0_cfi_flash_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_0_cfi_flash_uas_read,          --      .read
			uas_write            => mm_interconnect_0_cfi_flash_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_0_cfi_flash_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_0_cfi_flash_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_0_cfi_flash_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_0_cfi_flash_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_0_cfi_flash_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_0_cfi_flash_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_0_cfi_flash_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => cfi_flash_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_read_n_out       => cfi_flash_tcm_read_n_out,                      --      .read_n_out
			tcm_chipselect_n_out => cfi_flash_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => cfi_flash_tcm_request,                         --      .request
			tcm_grant            => cfi_flash_tcm_grant,                           --      .grant
			tcm_address_out      => cfi_flash_tcm_address_out,                     --      .address_out
			tcm_data_out         => cfi_flash_tcm_data_out,                        --      .data_out
			tcm_data_outen       => cfi_flash_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => cfi_flash_tcm_data_in                          --      .data_in
		);

	clock_crossing_io : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 9,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 32,
			RESPONSE_FIFO_DEPTH => 256,
			MASTER_SYNC_DEPTH   => 3,
			SLAVE_SYNC_DEPTH    => 3
		)
		port map (
			m0_clk           => altpll_c2_clk,                                        --   m0_clk.clk
			m0_reset         => rst_controller_003_reset_out_reset,                   -- m0_reset.reset
			s0_clk           => altpll_c0_clk,                                        --   s0_clk.clk
			s0_reset         => rst_controller_002_reset_out_reset,                   -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_clock_crossing_io_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_clock_crossing_io_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_clock_crossing_io_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_clock_crossing_io_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_clock_crossing_io_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_clock_crossing_io_s0_address,       --         .address
			s0_write         => mm_interconnect_0_clock_crossing_io_s0_write,         --         .write
			s0_read          => mm_interconnect_0_clock_crossing_io_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_clock_crossing_io_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_clock_crossing_io_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => clock_crossing_io_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => clock_crossing_io_m0_readdata,                        --         .readdata
			m0_readdatavalid => clock_crossing_io_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => clock_crossing_io_m0_burstcount,                      --         .burstcount
			m0_writedata     => clock_crossing_io_m0_writedata,                       --         .writedata
			m0_address       => clock_crossing_io_m0_address,                         --         .address
			m0_write         => clock_crossing_io_m0_write,                           --         .write
			m0_read          => clock_crossing_io_m0_read,                            --         .read
			m0_byteenable    => clock_crossing_io_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => clock_crossing_io_m0_debugaccess                      --         .debugaccess
		);

	cpu : component DE2_115_SD_CARD_NIOS_cpu
		port map (
			clk                                 => altpll_c0_clk,                                     --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	floatdata_output : component DE2_115_SD_CARD_NIOS_floatdata_output
		port map (
			clk        => altpll_c0_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_floatdata_output_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_floatdata_output_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_floatdata_output_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_floatdata_output_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_floatdata_output_s1_readdata,        --                    .readdata
			out_port   => floatdata_output_external_connection_export            -- external_connection.export
		);

	jtag_uart : component DE2_115_SD_CARD_NIOS_jtag_uart
		port map (
			clk            => altpll_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	key : component DE2_115_SD_CARD_NIOS_key
		port map (
			clk        => altpll_c0_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port    => key_external_connection_export            -- external_connection.export
		);

	ledg : component DE2_115_SD_CARD_NIOS_ledg
		port map (
			clk        => altpll_c0_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_ledg_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_ledg_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_ledg_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_ledg_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_ledg_s1_readdata,        --                    .readdata
			out_port   => ledg_external_connection_export            -- external_connection.export
		);

	ledr : component DE2_115_SD_CARD_NIOS_ledr
		port map (
			clk        => altpll_c0_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_ledr_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_ledr_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_ledr_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_ledr_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_ledr_s1_readdata,        --                    .readdata
			out_port   => ledr_external_connection_export            -- external_connection.export
		);

	onchip_memory2 : component DE2_115_SD_CARD_NIOS_onchip_memory2
		port map (
			clk        => altpll_c0_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,             --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	pixel_index : component DE2_115_SD_CARD_NIOS_pixel_index
		port map (
			clk        => altpll_c0_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_pixel_index_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pixel_index_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pixel_index_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pixel_index_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pixel_index_s1_readdata,        --                    .readdata
			out_port   => pixel_index_external_connection_export            -- external_connection.export
		);

	results_input : component DE2_115_SD_CARD_NIOS_results_input
		port map (
			clk      => altpll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => mm_interconnect_0_results_input_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_results_input_s1_readdata, --                    .readdata
			in_port  => results_input_external_connection_export     -- external_connection.export
		);

	sd_clk : component DE2_115_SD_CARD_NIOS_sd_clk
		port map (
			clk        => altpll_c0_clk,                                --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_sd_clk_s1_address,          --                  s1.address
			write_n    => mm_interconnect_1_sd_clk_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_1_sd_clk_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_1_sd_clk_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_1_sd_clk_s1_readdata,         --                    .readdata
			out_port   => sd_clk_external_connection_export             -- external_connection.export
		);

	sd_cmd : component DE2_115_SD_CARD_NIOS_sd_cmd
		port map (
			clk        => altpll_c0_clk,                                --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_sd_cmd_s1_address,          --                  s1.address
			write_n    => mm_interconnect_1_sd_cmd_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_1_sd_cmd_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_1_sd_cmd_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_1_sd_cmd_s1_readdata,         --                    .readdata
			bidir_port => sd_cmd_external_connection_export             -- external_connection.export
		);

	sd_dat : component DE2_115_SD_CARD_NIOS_sd_dat
		port map (
			clk        => altpll_c0_clk,                                --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_sd_dat_s1_address,          --                  s1.address
			write_n    => mm_interconnect_1_sd_dat_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_1_sd_dat_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_1_sd_dat_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_1_sd_dat_s1_readdata,         --                    .readdata
			bidir_port => sd_dat_external_connection_export             -- external_connection.export
		);

	sd_wp_n : component DE2_115_SD_CARD_NIOS_sd_wp_n
		port map (
			clk      => altpll_c0_clk,                                --                 clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_sd_wp_n_s1_address,         --                  s1.address
			readdata => mm_interconnect_1_sd_wp_n_s1_readdata,        --                    .readdata
			in_port  => sd_wp_n_external_connection_export            -- external_connection.export
		);

	sw : component DE2_115_SD_CARD_NIOS_sw
		port map (
			clk        => altpll_c0_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_sw_s1_address,          --                  s1.address
			write_n    => mm_interconnect_0_sw_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_0_sw_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_0_sw_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_0_sw_s1_readdata,         --                    .readdata
			in_port    => sw_external_connection_export             -- external_connection.export
		);

	sync_data : component DE2_115_SD_CARD_NIOS_sync_data
		port map (
			clk        => altpll_c0_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_sync_data_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sync_data_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sync_data_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sync_data_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sync_data_s1_readdata,        --                    .readdata
			out_port   => sync_data_external_connection_export            -- external_connection.export
		);

	timer : component DE2_115_SD_CARD_NIOS_timer
		port map (
			clk        => altpll_c0_clk,                                --   clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_1_timer_s1_address,           --    s1.address
			writedata  => mm_interconnect_1_timer_s1_writedata,         --      .writedata
			readdata   => mm_interconnect_1_timer_s1_readdata,          --      .readdata
			chipselect => mm_interconnect_1_timer_s1_chipselect,        --      .chipselect
			write_n    => mm_interconnect_1_timer_s1_write_ports_inv,   --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	tri_state_bridge_flash_bridge_0 : component DE2_115_SD_CARD_NIOS_tri_state_bridge_flash_bridge_0
		port map (
			clk                                   => altpll_c0_clk,                                                            --   clk.clk
			reset                                 => rst_controller_002_reset_out_reset,                                       -- reset.reset
			request                               => tri_state_flash_bridge_pinsharer_0_tcm_request,                           --   tcs.request
			grant                                 => tri_state_flash_bridge_pinsharer_0_tcm_grant,                             --      .grant
			tcs_address_to_the_cfi_flash          => tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out,      --      .address_to_the_cfi_flash_out
			tcs_tri_state_bridge_flash_data       => tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out,   --      .tri_state_bridge_flash_data_out
			tcs_tri_state_bridge_flash_data_outen => tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen, --      .tri_state_bridge_flash_data_outen
			tcs_tri_state_bridge_flash_data_in    => tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in,    --      .tri_state_bridge_flash_data_in
			tcs_write_n_to_the_cfi_flash          => tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out,      --      .write_n_to_the_cfi_flash_out
			tcs_select_n_to_the_cfi_flash         => tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out,     --      .select_n_to_the_cfi_flash_out
			tcs_read_n_to_the_cfi_flash           => tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out,       --      .read_n_to_the_cfi_flash_out
			address_to_the_cfi_flash              => tri_state_bridge_flash_bridge_0_out_address_to_the_cfi_flash,             --   out.address_to_the_cfi_flash
			tri_state_bridge_flash_data           => tri_state_bridge_flash_bridge_0_out_tri_state_bridge_flash_data,          --      .tri_state_bridge_flash_data
			write_n_to_the_cfi_flash              => tri_state_bridge_flash_bridge_0_out_write_n_to_the_cfi_flash,             --      .write_n_to_the_cfi_flash
			select_n_to_the_cfi_flash             => tri_state_bridge_flash_bridge_0_out_select_n_to_the_cfi_flash,            --      .select_n_to_the_cfi_flash
			read_n_to_the_cfi_flash               => tri_state_bridge_flash_bridge_0_out_read_n_to_the_cfi_flash               --      .read_n_to_the_cfi_flash
		);

	tri_state_flash_bridge_pinsharer_0 : component DE2_115_SD_CARD_NIOS_tri_state_flash_bridge_pinSharer_0
		port map (
			clk_clk                           => altpll_c0_clk,                                                            --   clk.clk
			reset_reset                       => rst_controller_002_reset_out_reset,                                       -- reset.reset
			request                           => tri_state_flash_bridge_pinsharer_0_tcm_request,                           --   tcm.request
			grant                             => tri_state_flash_bridge_pinsharer_0_tcm_grant,                             --      .grant
			address_to_the_cfi_flash          => tri_state_flash_bridge_pinsharer_0_tcm_address_to_the_cfi_flash_out,      --      .address_to_the_cfi_flash_out
			read_n_to_the_cfi_flash           => tri_state_flash_bridge_pinsharer_0_tcm_read_n_to_the_cfi_flash_out,       --      .read_n_to_the_cfi_flash_out
			write_n_to_the_cfi_flash          => tri_state_flash_bridge_pinsharer_0_tcm_write_n_to_the_cfi_flash_out,      --      .write_n_to_the_cfi_flash_out
			tri_state_bridge_flash_data       => tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_out,   --      .tri_state_bridge_flash_data_out
			tri_state_bridge_flash_data_in    => tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_in,    --      .tri_state_bridge_flash_data_in
			tri_state_bridge_flash_data_outen => tri_state_flash_bridge_pinsharer_0_tcm_tri_state_bridge_flash_data_outen, --      .tri_state_bridge_flash_data_outen
			select_n_to_the_cfi_flash         => tri_state_flash_bridge_pinsharer_0_tcm_select_n_to_the_cfi_flash_out,     --      .select_n_to_the_cfi_flash_out
			tcs0_request                      => cfi_flash_tcm_request,                                                    --  tcs0.request
			tcs0_grant                        => cfi_flash_tcm_grant,                                                      --      .grant
			tcs0_address_out                  => cfi_flash_tcm_address_out,                                                --      .address_out
			tcs0_read_n_out(0)                => cfi_flash_tcm_read_n_out,                                                 --      .read_n_out
			tcs0_write_n_out(0)               => cfi_flash_tcm_write_n_out,                                                --      .write_n_out
			tcs0_data_out                     => cfi_flash_tcm_data_out,                                                   --      .data_out
			tcs0_data_in                      => cfi_flash_tcm_data_in,                                                    --      .data_in
			tcs0_data_outen                   => cfi_flash_tcm_data_outen,                                                 --      .data_outen
			tcs0_chipselect_n_out(0)          => cfi_flash_tcm_chipselect_n_out                                            --      .chipselect_n_out
		);

	video_character_buffer_with_dma_0 : component DE2_115_SD_CARD_NIOS_video_character_buffer_with_dma_0
		port map (
			clk                  => video_pll_0_vga_clk_clk,                                                                    --                       clk.clk
			reset                => rst_controller_004_reset_out_reset,                                                         --                     reset.reset
			ctrl_address         => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address(0),   -- avalon_char_control_slave.address
			ctrl_byteenable      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable,   --                          .byteenable
			ctrl_chipselect      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect,   --                          .chipselect
			ctrl_read            => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read,         --                          .read
			ctrl_write           => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write,        --                          .write
			ctrl_writedata       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata,    --                          .writedata
			ctrl_readdata        => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata,     --                          .readdata
			buf_byteenable       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable(0), --  avalon_char_buffer_slave.byteenable
			buf_chipselect       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect,    --                          .chipselect
			buf_read             => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read,          --                          .read
			buf_write            => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write,         --                          .write
			buf_writedata        => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata,     --                          .writedata
			buf_readdata         => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata,      --                          .readdata
			buf_waitrequest      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest,   --                          .waitrequest
			buf_address          => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address,       --                          .address
			stream_ready         => video_character_buffer_with_dma_0_avalon_char_source_ready,                                 --        avalon_char_source.ready
			stream_startofpacket => video_character_buffer_with_dma_0_avalon_char_source_startofpacket,                         --                          .startofpacket
			stream_endofpacket   => video_character_buffer_with_dma_0_avalon_char_source_endofpacket,                           --                          .endofpacket
			stream_valid         => video_character_buffer_with_dma_0_avalon_char_source_valid,                                 --                          .valid
			stream_data          => video_character_buffer_with_dma_0_avalon_char_source_data                                   --                          .data
		);

	video_pll_0 : component DE2_115_SD_CARD_NIOS_video_pll_0
		port map (
			ref_clk_clk        => clk_50_clk_in_clk,                  --      ref_clk.clk
			ref_reset_reset    => rst_controller_005_reset_out_reset, --    ref_reset.reset
			vga_clk_clk        => video_pll_0_vga_clk_clk,            --      vga_clk.clk
			lcd_clk_clk        => open,                               --      lcd_clk.clk
			reset_source_reset => video_pll_0_reset_source_reset      -- reset_source.reset
		);

	video_vga_controller_0 : component DE2_115_SD_CARD_NIOS_video_vga_controller_0
		port map (
			clk           => video_pll_0_vga_clk_clk,                                            --                clk.clk
			reset         => rst_controller_004_reset_out_reset,                                 --              reset.reset
			data          => video_character_buffer_with_dma_0_avalon_char_source_data,          --    avalon_vga_sink.data
			startofpacket => video_character_buffer_with_dma_0_avalon_char_source_startofpacket, --                   .startofpacket
			endofpacket   => video_character_buffer_with_dma_0_avalon_char_source_endofpacket,   --                   .endofpacket
			valid         => video_character_buffer_with_dma_0_avalon_char_source_valid,         --                   .valid
			ready         => video_character_buffer_with_dma_0_avalon_char_source_ready,         --                   .ready
			VGA_CLK       => video_vga_controller_0_external_interface_CLK,                      -- external_interface.export
			VGA_HS        => video_vga_controller_0_external_interface_HS,                       --                   .export
			VGA_VS        => video_vga_controller_0_external_interface_VS,                       --                   .export
			VGA_BLANK     => video_vga_controller_0_external_interface_BLANK,                    --                   .export
			VGA_SYNC      => video_vga_controller_0_external_interface_SYNC,                     --                   .export
			VGA_R         => video_vga_controller_0_external_interface_R,                        --                   .export
			VGA_G         => video_vga_controller_0_external_interface_G,                        --                   .export
			VGA_B         => video_vga_controller_0_external_interface_B                         --                   .export
		);

	weight_index : component DE2_115_SD_CARD_NIOS_weight_index
		port map (
			clk        => altpll_c0_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_weight_index_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_weight_index_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_weight_index_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_weight_index_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_weight_index_s1_readdata,        --                    .readdata
			out_port   => weight_index_external_connection_export            -- external_connection.export
		);

	mm_interconnect_0 : component DE2_115_SD_CARD_NIOS_mm_interconnect_0
		port map (
			altpll_c0_clk                                                          => altpll_c0_clk,                                                                            --                                                     altpll_c0.clk
			clk_50_clk_clk                                                         => clk_50_clk_in_clk,                                                                        --                                                    clk_50_clk.clk
			video_pll_0_vga_clk_clk                                                => video_pll_0_vga_clk_clk,                                                                  --                                           video_pll_0_vga_clk.clk
			altpll_inclk_interface_reset_reset_bridge_in_reset_reset               => rst_controller_001_reset_out_reset,                                                       --            altpll_inclk_interface_reset_reset_bridge_in_reset.reset
			cpu_reset_reset_bridge_in_reset_reset                                  => rst_controller_002_reset_out_reset,                                                       --                               cpu_reset_reset_bridge_in_reset.reset
			onchip_memory2_reset1_reset_bridge_in_reset_reset                      => rst_controller_reset_out_reset,                                                           --                   onchip_memory2_reset1_reset_bridge_in_reset.reset
			video_character_buffer_with_dma_0_reset_reset_bridge_in_reset_reset    => rst_controller_004_reset_out_reset,                                                       -- video_character_buffer_with_dma_0_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                                => cpu_data_master_address,                                                                  --                                               cpu_data_master.address
			cpu_data_master_waitrequest                                            => cpu_data_master_waitrequest,                                                              --                                                              .waitrequest
			cpu_data_master_byteenable                                             => cpu_data_master_byteenable,                                                               --                                                              .byteenable
			cpu_data_master_read                                                   => cpu_data_master_read,                                                                     --                                                              .read
			cpu_data_master_readdata                                               => cpu_data_master_readdata,                                                                 --                                                              .readdata
			cpu_data_master_readdatavalid                                          => cpu_data_master_readdatavalid,                                                            --                                                              .readdatavalid
			cpu_data_master_write                                                  => cpu_data_master_write,                                                                    --                                                              .write
			cpu_data_master_writedata                                              => cpu_data_master_writedata,                                                                --                                                              .writedata
			cpu_data_master_debugaccess                                            => cpu_data_master_debugaccess,                                                              --                                                              .debugaccess
			cpu_instruction_master_address                                         => cpu_instruction_master_address,                                                           --                                        cpu_instruction_master.address
			cpu_instruction_master_waitrequest                                     => cpu_instruction_master_waitrequest,                                                       --                                                              .waitrequest
			cpu_instruction_master_read                                            => cpu_instruction_master_read,                                                              --                                                              .read
			cpu_instruction_master_readdata                                        => cpu_instruction_master_readdata,                                                          --                                                              .readdata
			cpu_instruction_master_readdatavalid                                   => cpu_instruction_master_readdatavalid,                                                     --                                                              .readdatavalid
			activations_index_s1_address                                           => mm_interconnect_0_activations_index_s1_address,                                           --                                          activations_index_s1.address
			activations_index_s1_write                                             => mm_interconnect_0_activations_index_s1_write,                                             --                                                              .write
			activations_index_s1_readdata                                          => mm_interconnect_0_activations_index_s1_readdata,                                          --                                                              .readdata
			activations_index_s1_writedata                                         => mm_interconnect_0_activations_index_s1_writedata,                                         --                                                              .writedata
			activations_index_s1_chipselect                                        => mm_interconnect_0_activations_index_s1_chipselect,                                        --                                                              .chipselect
			altpll_pll_slave_address                                               => mm_interconnect_0_altpll_pll_slave_address,                                               --                                              altpll_pll_slave.address
			altpll_pll_slave_write                                                 => mm_interconnect_0_altpll_pll_slave_write,                                                 --                                                              .write
			altpll_pll_slave_read                                                  => mm_interconnect_0_altpll_pll_slave_read,                                                  --                                                              .read
			altpll_pll_slave_readdata                                              => mm_interconnect_0_altpll_pll_slave_readdata,                                              --                                                              .readdata
			altpll_pll_slave_writedata                                             => mm_interconnect_0_altpll_pll_slave_writedata,                                             --                                                              .writedata
			cfi_flash_uas_address                                                  => mm_interconnect_0_cfi_flash_uas_address,                                                  --                                                 cfi_flash_uas.address
			cfi_flash_uas_write                                                    => mm_interconnect_0_cfi_flash_uas_write,                                                    --                                                              .write
			cfi_flash_uas_read                                                     => mm_interconnect_0_cfi_flash_uas_read,                                                     --                                                              .read
			cfi_flash_uas_readdata                                                 => mm_interconnect_0_cfi_flash_uas_readdata,                                                 --                                                              .readdata
			cfi_flash_uas_writedata                                                => mm_interconnect_0_cfi_flash_uas_writedata,                                                --                                                              .writedata
			cfi_flash_uas_burstcount                                               => mm_interconnect_0_cfi_flash_uas_burstcount,                                               --                                                              .burstcount
			cfi_flash_uas_byteenable                                               => mm_interconnect_0_cfi_flash_uas_byteenable,                                               --                                                              .byteenable
			cfi_flash_uas_readdatavalid                                            => mm_interconnect_0_cfi_flash_uas_readdatavalid,                                            --                                                              .readdatavalid
			cfi_flash_uas_waitrequest                                              => mm_interconnect_0_cfi_flash_uas_waitrequest,                                              --                                                              .waitrequest
			cfi_flash_uas_lock                                                     => mm_interconnect_0_cfi_flash_uas_lock,                                                     --                                                              .lock
			cfi_flash_uas_debugaccess                                              => mm_interconnect_0_cfi_flash_uas_debugaccess,                                              --                                                              .debugaccess
			clock_crossing_io_s0_address                                           => mm_interconnect_0_clock_crossing_io_s0_address,                                           --                                          clock_crossing_io_s0.address
			clock_crossing_io_s0_write                                             => mm_interconnect_0_clock_crossing_io_s0_write,                                             --                                                              .write
			clock_crossing_io_s0_read                                              => mm_interconnect_0_clock_crossing_io_s0_read,                                              --                                                              .read
			clock_crossing_io_s0_readdata                                          => mm_interconnect_0_clock_crossing_io_s0_readdata,                                          --                                                              .readdata
			clock_crossing_io_s0_writedata                                         => mm_interconnect_0_clock_crossing_io_s0_writedata,                                         --                                                              .writedata
			clock_crossing_io_s0_burstcount                                        => mm_interconnect_0_clock_crossing_io_s0_burstcount,                                        --                                                              .burstcount
			clock_crossing_io_s0_byteenable                                        => mm_interconnect_0_clock_crossing_io_s0_byteenable,                                        --                                                              .byteenable
			clock_crossing_io_s0_readdatavalid                                     => mm_interconnect_0_clock_crossing_io_s0_readdatavalid,                                     --                                                              .readdatavalid
			clock_crossing_io_s0_waitrequest                                       => mm_interconnect_0_clock_crossing_io_s0_waitrequest,                                       --                                                              .waitrequest
			clock_crossing_io_s0_debugaccess                                       => mm_interconnect_0_clock_crossing_io_s0_debugaccess,                                       --                                                              .debugaccess
			cpu_debug_mem_slave_address                                            => mm_interconnect_0_cpu_debug_mem_slave_address,                                            --                                           cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                              => mm_interconnect_0_cpu_debug_mem_slave_write,                                              --                                                              .write
			cpu_debug_mem_slave_read                                               => mm_interconnect_0_cpu_debug_mem_slave_read,                                               --                                                              .read
			cpu_debug_mem_slave_readdata                                           => mm_interconnect_0_cpu_debug_mem_slave_readdata,                                           --                                                              .readdata
			cpu_debug_mem_slave_writedata                                          => mm_interconnect_0_cpu_debug_mem_slave_writedata,                                          --                                                              .writedata
			cpu_debug_mem_slave_byteenable                                         => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                                         --                                                              .byteenable
			cpu_debug_mem_slave_waitrequest                                        => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                                        --                                                              .waitrequest
			cpu_debug_mem_slave_debugaccess                                        => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                                        --                                                              .debugaccess
			floatdata_output_s1_address                                            => mm_interconnect_0_floatdata_output_s1_address,                                            --                                           floatdata_output_s1.address
			floatdata_output_s1_write                                              => mm_interconnect_0_floatdata_output_s1_write,                                              --                                                              .write
			floatdata_output_s1_readdata                                           => mm_interconnect_0_floatdata_output_s1_readdata,                                           --                                                              .readdata
			floatdata_output_s1_writedata                                          => mm_interconnect_0_floatdata_output_s1_writedata,                                          --                                                              .writedata
			floatdata_output_s1_chipselect                                         => mm_interconnect_0_floatdata_output_s1_chipselect,                                         --                                                              .chipselect
			jtag_uart_avalon_jtag_slave_address                                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,                                    --                                   jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                                      --                                                              .write
			jtag_uart_avalon_jtag_slave_read                                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                                       --                                                              .read
			jtag_uart_avalon_jtag_slave_readdata                                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,                                   --                                                              .readdata
			jtag_uart_avalon_jtag_slave_writedata                                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,                                  --                                                              .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,                                --                                                              .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,                                 --                                                              .chipselect
			key_s1_address                                                         => mm_interconnect_0_key_s1_address,                                                         --                                                        key_s1.address
			key_s1_write                                                           => mm_interconnect_0_key_s1_write,                                                           --                                                              .write
			key_s1_readdata                                                        => mm_interconnect_0_key_s1_readdata,                                                        --                                                              .readdata
			key_s1_writedata                                                       => mm_interconnect_0_key_s1_writedata,                                                       --                                                              .writedata
			key_s1_chipselect                                                      => mm_interconnect_0_key_s1_chipselect,                                                      --                                                              .chipselect
			ledg_s1_address                                                        => mm_interconnect_0_ledg_s1_address,                                                        --                                                       ledg_s1.address
			ledg_s1_write                                                          => mm_interconnect_0_ledg_s1_write,                                                          --                                                              .write
			ledg_s1_readdata                                                       => mm_interconnect_0_ledg_s1_readdata,                                                       --                                                              .readdata
			ledg_s1_writedata                                                      => mm_interconnect_0_ledg_s1_writedata,                                                      --                                                              .writedata
			ledg_s1_chipselect                                                     => mm_interconnect_0_ledg_s1_chipselect,                                                     --                                                              .chipselect
			ledr_s1_address                                                        => mm_interconnect_0_ledr_s1_address,                                                        --                                                       ledr_s1.address
			ledr_s1_write                                                          => mm_interconnect_0_ledr_s1_write,                                                          --                                                              .write
			ledr_s1_readdata                                                       => mm_interconnect_0_ledr_s1_readdata,                                                       --                                                              .readdata
			ledr_s1_writedata                                                      => mm_interconnect_0_ledr_s1_writedata,                                                      --                                                              .writedata
			ledr_s1_chipselect                                                     => mm_interconnect_0_ledr_s1_chipselect,                                                     --                                                              .chipselect
			onchip_memory2_s1_address                                              => mm_interconnect_0_onchip_memory2_s1_address,                                              --                                             onchip_memory2_s1.address
			onchip_memory2_s1_write                                                => mm_interconnect_0_onchip_memory2_s1_write,                                                --                                                              .write
			onchip_memory2_s1_readdata                                             => mm_interconnect_0_onchip_memory2_s1_readdata,                                             --                                                              .readdata
			onchip_memory2_s1_writedata                                            => mm_interconnect_0_onchip_memory2_s1_writedata,                                            --                                                              .writedata
			onchip_memory2_s1_byteenable                                           => mm_interconnect_0_onchip_memory2_s1_byteenable,                                           --                                                              .byteenable
			onchip_memory2_s1_chipselect                                           => mm_interconnect_0_onchip_memory2_s1_chipselect,                                           --                                                              .chipselect
			onchip_memory2_s1_clken                                                => mm_interconnect_0_onchip_memory2_s1_clken,                                                --                                                              .clken
			pixel_index_s1_address                                                 => mm_interconnect_0_pixel_index_s1_address,                                                 --                                                pixel_index_s1.address
			pixel_index_s1_write                                                   => mm_interconnect_0_pixel_index_s1_write,                                                   --                                                              .write
			pixel_index_s1_readdata                                                => mm_interconnect_0_pixel_index_s1_readdata,                                                --                                                              .readdata
			pixel_index_s1_writedata                                               => mm_interconnect_0_pixel_index_s1_writedata,                                               --                                                              .writedata
			pixel_index_s1_chipselect                                              => mm_interconnect_0_pixel_index_s1_chipselect,                                              --                                                              .chipselect
			results_input_s1_address                                               => mm_interconnect_0_results_input_s1_address,                                               --                                              results_input_s1.address
			results_input_s1_readdata                                              => mm_interconnect_0_results_input_s1_readdata,                                              --                                                              .readdata
			sw_s1_address                                                          => mm_interconnect_0_sw_s1_address,                                                          --                                                         sw_s1.address
			sw_s1_write                                                            => mm_interconnect_0_sw_s1_write,                                                            --                                                              .write
			sw_s1_readdata                                                         => mm_interconnect_0_sw_s1_readdata,                                                         --                                                              .readdata
			sw_s1_writedata                                                        => mm_interconnect_0_sw_s1_writedata,                                                        --                                                              .writedata
			sw_s1_chipselect                                                       => mm_interconnect_0_sw_s1_chipselect,                                                       --                                                              .chipselect
			sync_data_s1_address                                                   => mm_interconnect_0_sync_data_s1_address,                                                   --                                                  sync_data_s1.address
			sync_data_s1_write                                                     => mm_interconnect_0_sync_data_s1_write,                                                     --                                                              .write
			sync_data_s1_readdata                                                  => mm_interconnect_0_sync_data_s1_readdata,                                                  --                                                              .readdata
			sync_data_s1_writedata                                                 => mm_interconnect_0_sync_data_s1_writedata,                                                 --                                                              .writedata
			sync_data_s1_chipselect                                                => mm_interconnect_0_sync_data_s1_chipselect,                                                --                                                              .chipselect
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address,     --    video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write,       --                                                              .write
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read,        --                                                              .read
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata,    --                                                              .readdata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata,   --                                                              .writedata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable,  --                                                              .byteenable
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest, --                                                              .waitrequest
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect,  --                                                              .chipselect
			video_character_buffer_with_dma_0_avalon_char_control_slave_address    => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address,    --   video_character_buffer_with_dma_0_avalon_char_control_slave.address
			video_character_buffer_with_dma_0_avalon_char_control_slave_write      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write,      --                                                              .write
			video_character_buffer_with_dma_0_avalon_char_control_slave_read       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read,       --                                                              .read
			video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata,   --                                                              .readdata
			video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata,  --                                                              .writedata
			video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable, --                                                              .byteenable
			video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect, --                                                              .chipselect
			weight_index_s1_address                                                => mm_interconnect_0_weight_index_s1_address,                                                --                                               weight_index_s1.address
			weight_index_s1_write                                                  => mm_interconnect_0_weight_index_s1_write,                                                  --                                                              .write
			weight_index_s1_readdata                                               => mm_interconnect_0_weight_index_s1_readdata,                                               --                                                              .readdata
			weight_index_s1_writedata                                              => mm_interconnect_0_weight_index_s1_writedata,                                              --                                                              .writedata
			weight_index_s1_chipselect                                             => mm_interconnect_0_weight_index_s1_chipselect                                              --                                                              .chipselect
		);

	mm_interconnect_1 : component DE2_115_SD_CARD_NIOS_mm_interconnect_1
		port map (
			altpll_c0_clk                                          => altpll_c0_clk,                          --                                        altpll_c0.clk
			altpll_c2_clk                                          => altpll_c2_clk,                          --                                        altpll_c2.clk
			clock_crossing_io_m0_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,     -- clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
			sd_clk_reset_reset_bridge_in_reset_reset               => rst_controller_002_reset_out_reset,     --               sd_clk_reset_reset_bridge_in_reset.reset
			clock_crossing_io_m0_address                           => clock_crossing_io_m0_address,           --                             clock_crossing_io_m0.address
			clock_crossing_io_m0_waitrequest                       => clock_crossing_io_m0_waitrequest,       --                                                 .waitrequest
			clock_crossing_io_m0_burstcount                        => clock_crossing_io_m0_burstcount,        --                                                 .burstcount
			clock_crossing_io_m0_byteenable                        => clock_crossing_io_m0_byteenable,        --                                                 .byteenable
			clock_crossing_io_m0_read                              => clock_crossing_io_m0_read,              --                                                 .read
			clock_crossing_io_m0_readdata                          => clock_crossing_io_m0_readdata,          --                                                 .readdata
			clock_crossing_io_m0_readdatavalid                     => clock_crossing_io_m0_readdatavalid,     --                                                 .readdatavalid
			clock_crossing_io_m0_write                             => clock_crossing_io_m0_write,             --                                                 .write
			clock_crossing_io_m0_writedata                         => clock_crossing_io_m0_writedata,         --                                                 .writedata
			clock_crossing_io_m0_debugaccess                       => clock_crossing_io_m0_debugaccess,       --                                                 .debugaccess
			sd_clk_s1_address                                      => mm_interconnect_1_sd_clk_s1_address,    --                                        sd_clk_s1.address
			sd_clk_s1_write                                        => mm_interconnect_1_sd_clk_s1_write,      --                                                 .write
			sd_clk_s1_readdata                                     => mm_interconnect_1_sd_clk_s1_readdata,   --                                                 .readdata
			sd_clk_s1_writedata                                    => mm_interconnect_1_sd_clk_s1_writedata,  --                                                 .writedata
			sd_clk_s1_chipselect                                   => mm_interconnect_1_sd_clk_s1_chipselect, --                                                 .chipselect
			sd_cmd_s1_address                                      => mm_interconnect_1_sd_cmd_s1_address,    --                                        sd_cmd_s1.address
			sd_cmd_s1_write                                        => mm_interconnect_1_sd_cmd_s1_write,      --                                                 .write
			sd_cmd_s1_readdata                                     => mm_interconnect_1_sd_cmd_s1_readdata,   --                                                 .readdata
			sd_cmd_s1_writedata                                    => mm_interconnect_1_sd_cmd_s1_writedata,  --                                                 .writedata
			sd_cmd_s1_chipselect                                   => mm_interconnect_1_sd_cmd_s1_chipselect, --                                                 .chipselect
			sd_dat_s1_address                                      => mm_interconnect_1_sd_dat_s1_address,    --                                        sd_dat_s1.address
			sd_dat_s1_write                                        => mm_interconnect_1_sd_dat_s1_write,      --                                                 .write
			sd_dat_s1_readdata                                     => mm_interconnect_1_sd_dat_s1_readdata,   --                                                 .readdata
			sd_dat_s1_writedata                                    => mm_interconnect_1_sd_dat_s1_writedata,  --                                                 .writedata
			sd_dat_s1_chipselect                                   => mm_interconnect_1_sd_dat_s1_chipselect, --                                                 .chipselect
			sd_wp_n_s1_address                                     => mm_interconnect_1_sd_wp_n_s1_address,   --                                       sd_wp_n_s1.address
			sd_wp_n_s1_readdata                                    => mm_interconnect_1_sd_wp_n_s1_readdata,  --                                                 .readdata
			timer_s1_address                                       => mm_interconnect_1_timer_s1_address,     --                                         timer_s1.address
			timer_s1_write                                         => mm_interconnect_1_timer_s1_write,       --                                                 .write
			timer_s1_readdata                                      => mm_interconnect_1_timer_s1_readdata,    --                                                 .readdata
			timer_s1_writedata                                     => mm_interconnect_1_timer_s1_writedata,   --                                                 .writedata
			timer_s1_chipselect                                    => mm_interconnect_1_timer_s1_chipselect   --                                                 .chipselect
		);

	irq_mapper : component DE2_115_SD_CARD_NIOS_irq_mapper
		port map (
			clk           => altpll_c0_clk,                      --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	rst_controller : component de2_115_sd_card_nios_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_c0_clk,                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component de2_115_sd_card_nios_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_50_clk_in_clk,                  --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component de2_115_sd_card_nios_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,          -- reset_in1.reset
			clk            => altpll_c0_clk,                          --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component de2_115_sd_card_nios_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => altpll_c2_clk,                      --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component de2_115_sd_card_nios_rst_controller_004
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => video_pll_0_reset_source_reset,     -- reset_in0.reset
			clk            => video_pll_0_vga_clk_clk,            --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_005 : component de2_115_sd_card_nios_rst_controller_004
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_50_clk_in_clk,                  --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_ledr_s1_write_ports_inv <= not mm_interconnect_0_ledr_s1_write;

	mm_interconnect_0_ledg_s1_write_ports_inv <= not mm_interconnect_0_ledg_s1_write;

	mm_interconnect_0_sw_s1_write_ports_inv <= not mm_interconnect_0_sw_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	mm_interconnect_0_floatdata_output_s1_write_ports_inv <= not mm_interconnect_0_floatdata_output_s1_write;

	mm_interconnect_0_sync_data_s1_write_ports_inv <= not mm_interconnect_0_sync_data_s1_write;

	mm_interconnect_0_pixel_index_s1_write_ports_inv <= not mm_interconnect_0_pixel_index_s1_write;

	mm_interconnect_0_weight_index_s1_write_ports_inv <= not mm_interconnect_0_weight_index_s1_write;

	mm_interconnect_0_activations_index_s1_write_ports_inv <= not mm_interconnect_0_activations_index_s1_write;

	mm_interconnect_1_sd_clk_s1_write_ports_inv <= not mm_interconnect_1_sd_clk_s1_write;

	mm_interconnect_1_sd_cmd_s1_write_ports_inv <= not mm_interconnect_1_sd_cmd_s1_write;

	mm_interconnect_1_sd_dat_s1_write_ports_inv <= not mm_interconnect_1_sd_dat_s1_write;

	mm_interconnect_1_timer_s1_write_ports_inv <= not mm_interconnect_1_timer_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	c0_out_clk_clk <= altpll_c0_clk;

	c2_out_clk_clk <= altpll_c2_clk;

end architecture rtl; -- of DE2_115_SD_CARD_NIOS
